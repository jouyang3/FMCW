library verilog;
use verilog.vl_types.all;
entity tb_memory is
end tb_memory;
