library verilog;
use verilog.vl_types.all;
entity tb_radar_top is
end tb_radar_top;
