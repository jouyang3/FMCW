library verilog;
use verilog.vl_types.all;
entity pll_testbench is
end pll_testbench;
