library verilog;
use verilog.vl_types.all;
entity tb_window is
end tb_window;
