library verilog;
use verilog.vl_types.all;
entity tb_magnitude is
end tb_magnitude;
