library verilog;
use verilog.vl_types.all;
entity dft_testbench is
end dft_testbench;
