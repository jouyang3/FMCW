library verilog;
use verilog.vl_types.all;
entity tb_FFT_Mag is
end tb_FFT_Mag;
