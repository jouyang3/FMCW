library verilog;
use verilog.vl_types.all;
entity tb_avg_filter is
end tb_avg_filter;
